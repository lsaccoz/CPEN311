module card7seg (card, seg7);

input [3:0] card;
output [6:0] seg7;
	
   // Your code for card7seg goes here. You can basically take the code directly
   // from your solution to Phase 2 (but notice that the inputs and outputs have
   // different names here).  Recall from Phase 2 that this is a purely 
   // combinational block.  

endmodule
