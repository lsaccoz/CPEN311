module statemachine ( slow_clock, resetb,
                      dscore, pscore, pcard3,
                      load_pcard1, load_pcard2,load_pcard3,
                      load_dcard1, load_dcard2, load_dcard3,
                      player_win_light, dealer_win_light);
							 
input slow_clock, resetb;
input [3:0] dscore, pscore, pcard3;
output reg load_pcard1, load_pcard2, load_pcard3;
output reg load_dcard1, load_dcard2, load_dcard3;
output reg player_win_light, dealer_win_light;


// The code describing your state machine will go here.  Remember that
// a state machine consists of next state logic, output logic, and the 
// registers that hold the state.  You will want to review your notes from
// CPEN 211 or equivalent if you have forgotten how to write a state machine.

wire [4:0] present_state;
reg [4:0] next_state;

DFF_5 state(.clk(slow_clock), .in(next_state), .out(present_state), .resetb(resetb));

	always @(*) begin
		case (present_state)
			5'd0: {next_state, load_dcard1, load_dcard2, load_dcard3, load_pcard1, load_pcard2, load_pcard3, player_win_light, dealer_win_light} = {5'd1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0};
			5'd1: {next_state, load_dcard1, load_dcard2, load_dcard3, load_pcard1, load_pcard2, load_pcard3, player_win_light, dealer_win_light} = {5'd2,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
			5'd2: {next_state, load_dcard1, load_dcard2, load_dcard3, load_pcard1, load_pcard2, load_pcard3, player_win_light, dealer_win_light} = {5'd3,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0};
			5'd3: {next_state, load_dcard1, load_dcard2, load_dcard3, load_pcard1, load_pcard2, load_pcard3, player_win_light, dealer_win_light} = {5'd4,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
			5'd4: begin
				{load_dcard1, load_dcard2, load_pcard1, load_pcard2, player_win_light, dealer_win_light} = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
				
				if(pscore>=4'd8 || dscore>=4'd8) begin
					next_state=5'd5;
					load_dcard3=1'b0;
					load_pcard3=1'b0;
				end
				else if((pscore==4'd6 || pscore==4'd7) && dscore<=4'd5) begin
					next_state=5'd5;
					load_dcard3=1'b1;
					load_pcard3=1'b0;
				end
				else if(pscore<=4'd5) begin
					next_state=5'd6;
					load_dcard3=1'b0;
					load_pcard3=1'b1;
				end
				else begin 
					next_state=5'd5;
					load_dcard3=1'b0;
					load_pcard3=1'b0;
				end
			end
			5'd5: begin 
				{next_state, load_dcard1, load_dcard2, load_dcard3, load_pcard1, load_pcard2, load_pcard3} = {5'd5,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
				if(pscore<dscore)
					{player_win_light,dealer_win_light} = 2'b01;
				else if (pscore>dscore)
					{player_win_light,dealer_win_light} = 2'b10;
				else
					{player_win_light,dealer_win_light} = 2'b11;
			end
			5'd6: begin 
				{next_state, load_dcard1, load_dcard2, load_pcard1, load_pcard2, load_pcard3, player_win_light, dealer_win_light} = {5'd5,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
				if(pcard3==4'd9&&dscore<=4'd3)
					load_dcard3=1'b1;
				else if(pcard3==4'd8&&dscore<=4'd2)
					load_dcard3=1'b1;
				else if(dscore<=((pcard3/2)+3) && pcard3<=4'd7)
					load_dcard3=1'b1;
				else
					load_dcard3=1'b0;
			end
			default:{next_state, load_dcard1, load_dcard2, load_dcard3, load_pcard1, load_pcard2, load_pcard3, player_win_light, dealer_win_light} = {5'd0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
		endcase
	end
endmodule

module DFF_5(clk, in, out, resetb) ;
	input clk, resetb;
	input [4:0] in;
	output reg [4:0] out;
	
	always @(posedge clk or negedge resetb) begin
		if(~resetb) begin
			out<=4'd0;
		end
		else
			out = in ;
	end
endmodule
			